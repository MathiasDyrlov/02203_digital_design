`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 11.09.2025 08:28:27
// Design Name: 
// Module Name: Talker_FSM
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module Talker_FSM(
    input clk,
    input reset,
    input start,
    input ack_sync,
    output ready,
    output req_out
    );
endmodule
